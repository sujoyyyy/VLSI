magic
tech scmos
timestamp 1596733371
<< nwell >>
rect -15 2 16 15
<< polysilicon >>
rect -1 13 1 17
rect -1 -5 1 4
rect -7 -8 1 -5
rect -1 -19 1 -8
rect -1 -30 1 -28
<< ndiffusion >>
rect -12 -20 -1 -19
rect -12 -24 -8 -20
rect -4 -24 -1 -20
rect -12 -28 -1 -24
rect 1 -22 13 -19
rect 1 -26 5 -22
rect 9 -26 13 -22
rect 1 -28 13 -26
<< pdiffusion >>
rect -12 9 -1 13
rect -12 5 -9 9
rect -5 5 -1 9
rect -12 4 -1 5
rect 1 11 13 13
rect 1 7 5 11
rect 9 7 13 11
rect 1 4 13 7
<< metal1 >>
rect -10 22 -6 26
rect -2 22 1 26
rect 5 22 9 26
rect -9 9 -5 22
rect 5 -5 9 7
rect 5 -8 14 -5
rect -8 -37 -4 -24
rect 5 -22 9 -8
rect -9 -41 -5 -37
rect -1 -41 3 -37
rect 7 -41 11 -37
<< ntransistor >>
rect -1 -28 1 -19
<< ptransistor >>
rect -1 4 1 13
<< ndcontact >>
rect -8 -24 -4 -20
rect 5 -26 9 -22
<< pdcontact >>
rect -9 5 -5 9
rect 5 7 9 11
<< emittercontact >>
rect 1 22 5 26
<< psubstratepcontact >>
rect -13 -41 -9 -37
rect -5 -41 -1 -37
rect 3 -41 7 -37
rect 11 -41 15 -37
<< nsubstratencontact >>
rect -14 22 -10 26
rect -6 22 -2 26
rect 9 22 13 26
<< labels >>
rlabel metal1 -9 24 -9 24 5 vdd
rlabel metal1 -7 -33 -7 -33 1 gnd
rlabel polysilicon -5 -7 -5 -7 1 vin
rlabel metal1 11 -7 11 -7 7 vout
<< end >>

module smallCircle(
    input Gi,
    output Ci
);
	
	buf buf0 (Ci, Gi);
	
endmodule

magic
tech scmos
timestamp 1596976683
<< nwell >>
rect -6 0 68 17
<< polysilicon >>
rect 6 7 8 9
rect 19 7 21 9
rect 29 7 31 9
rect 50 7 52 9
rect 6 -21 8 3
rect 19 -21 21 3
rect 29 -21 31 3
rect 50 -21 52 3
rect 6 -29 8 -26
rect 19 -29 21 -26
rect 29 -29 31 -26
rect 50 -29 52 -26
<< ndiffusion >>
rect 0 -26 1 -21
rect 5 -26 6 -21
rect 8 -26 19 -21
rect 21 -26 29 -21
rect 31 -26 33 -21
rect 37 -26 39 -21
rect 43 -26 44 -21
rect 48 -26 50 -21
rect 52 -26 56 -21
rect 60 -26 63 -21
<< pdiffusion >>
rect -1 3 0 7
rect 4 3 6 7
rect 8 3 13 7
rect 17 3 19 7
rect 21 3 22 7
rect 26 3 29 7
rect 31 3 33 7
rect 43 3 44 7
rect 48 3 50 7
rect 52 3 56 7
rect 60 3 63 7
<< metal1 >>
rect -5 13 -4 17
rect 0 7 4 17
rect 8 13 18 17
rect 22 7 26 17
rect 30 13 41 17
rect 45 13 49 17
rect 53 13 58 17
rect 62 13 65 17
rect 44 7 48 13
rect 13 -2 17 3
rect 33 -2 37 3
rect 13 -7 45 -2
rect 56 -5 60 3
rect -2 -15 2 -11
rect 11 -15 15 -11
rect 22 -15 25 -11
rect 33 -21 37 -7
rect 56 -9 66 -5
rect 56 -21 60 -9
rect 1 -36 5 -26
rect 44 -31 48 -26
rect 9 -36 15 -31
rect 19 -36 25 -31
rect 29 -36 40 -31
rect 44 -36 49 -31
rect 53 -36 58 -31
rect 62 -36 66 -31
<< ntransistor >>
rect 6 -26 8 -21
rect 19 -26 21 -21
rect 29 -26 31 -21
rect 50 -26 52 -21
<< ptransistor >>
rect 6 3 8 7
rect 19 3 21 7
rect 29 3 31 7
rect 50 3 52 7
<< polycontact >>
rect 2 -15 6 -11
rect 15 -15 19 -11
rect 25 -15 29 -11
rect 45 -7 50 -2
<< ndcontact >>
rect 1 -26 5 -21
rect 33 -26 37 -21
rect 44 -26 48 -21
rect 56 -26 60 -21
<< pdcontact >>
rect 0 3 4 7
rect 13 3 17 7
rect 22 3 26 7
rect 33 3 37 7
rect 44 3 48 7
rect 56 3 60 7
<< psubstratepcontact >>
rect -3 -36 1 -31
rect 5 -36 9 -31
rect 15 -36 19 -31
rect 25 -36 29 -31
rect 40 -36 44 -31
rect 49 -36 53 -31
rect 58 -36 62 -31
<< nsubstratencontact >>
rect -4 13 0 17
rect 4 13 8 17
rect 18 13 22 17
rect 26 13 30 17
rect 41 13 45 17
rect 49 13 53 17
rect 58 13 62 17
<< labels >>
rlabel metal1 12 -34 12 -34 1 gnd
rlabel metal1 36 -7 36 -2 1 out
rlabel metal1 66 -9 66 -5 7 Y
rlabel metal1 13 15 13 15 5 vdd
rlabel metal1 -1 -14 -1 -14 3 a
rlabel metal1 12 -14 12 -14 1 b
rlabel metal1 23 -14 23 -14 1 c
<< end >>
